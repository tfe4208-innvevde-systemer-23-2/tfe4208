
module DE2_115_SOPC (
	clk_clk,
	pwm_0_conduit_end_pwm,
	pwm_1_conduit_end_pwm,
	reset_reset_n);	

	input		clk_clk;
	output		pwm_0_conduit_end_pwm;
	output		pwm_1_conduit_end_pwm;
	input		reset_reset_n;
endmodule
