// Copyright

module Correlation_test;

endmodule;