
module DE2_115_SOPC (
	clk_clk,
	reset_reset_n,
	pwm_1_conduit_end_pwm,
	pwm_0_conduit_end_pwm);	

	input		clk_clk;
	input		reset_reset_n;
	output		pwm_1_conduit_end_pwm;
	output		pwm_0_conduit_end_pwm;
endmodule
