// Copyright

module Peak #(
    parameter MAX_LAGS                  = 17;
    parameter NUM_XCORRS                = 6;
) (
    input  logic                                    clk;
    input  logic                                    rst;
    
);

// Need edge detector???

endmodule