// Copyright

module CpuPeripheral_test;

endmodule;