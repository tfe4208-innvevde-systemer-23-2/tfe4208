// Copyright

module Peak_test;

endmodule;