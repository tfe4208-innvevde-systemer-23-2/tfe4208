// Copyright

module Mem_test;

endmodule;